magic
tech scmos
timestamp 1695278485
<< nwell >>
rect -4 6 17 18
<< polysilicon >>
rect 8 15 10 17
rect 8 5 10 9
rect 7 1 10 5
rect 8 -1 10 1
rect 8 -9 10 -7
<< ndiffusion >>
rect 3 -2 8 -1
rect 7 -6 8 -2
rect 3 -7 8 -6
rect 10 -2 15 -1
rect 10 -6 11 -2
rect 10 -7 15 -6
<< pdiffusion >>
rect 3 14 8 15
rect 7 10 8 14
rect 3 9 8 10
rect 10 14 15 15
rect 10 10 11 14
rect 10 9 15 10
<< metal1 >>
rect -3 21 15 25
rect 3 14 7 21
rect -3 1 3 5
rect 11 -2 15 10
rect 3 -13 7 -6
rect -3 -17 15 -13
<< ntransistor >>
rect 8 -7 10 -1
<< ptransistor >>
rect 8 9 10 15
<< polycontact >>
rect 3 1 7 5
<< ndcontact >>
rect 3 -6 7 -2
rect 11 -6 15 -2
<< pdcontact >>
rect 3 10 7 14
rect 11 10 15 14
<< psubstratepcontact >>
rect -1 -6 3 -2
<< nsubstratencontact >>
rect -1 10 3 14
<< labels >>
rlabel metal1 1 22 1 22 4 vdd
rlabel metal1 -1 3 -1 3 3 in
rlabel metal1 13 3 13 3 7 out
rlabel metal1 5 -15 5 -15 1 gnd
<< end >>
