magic
tech scmos
timestamp 1699438773
<< nwell >>
rect -18 -15 12 -4
<< polysilicon >>
rect -3 21 -1 23
rect -3 12 -1 15
rect -3 -7 -1 -3
rect -3 -15 -1 -13
<< ndiffusion >>
rect -10 20 -3 21
rect -10 16 -9 20
rect -5 16 -3 20
rect -10 15 -3 16
rect -1 20 7 21
rect -1 16 2 20
rect 6 16 7 20
rect -1 15 7 16
<< pdiffusion >>
rect -10 -8 -3 -7
rect -10 -12 -9 -8
rect -5 -12 -3 -8
rect -10 -13 -3 -12
rect -1 -8 7 -7
rect -1 -12 2 -8
rect 6 -12 7 -8
rect -1 -13 7 -12
<< metal1 >>
rect -33 24 -9 28
rect -9 20 -5 24
rect -33 16 -20 20
rect -33 8 -5 12
rect 2 8 6 16
rect 2 4 14 8
rect -33 -3 -5 1
rect 2 -8 6 4
rect -33 -12 -18 -8
rect -9 -17 -5 -12
<< metal2 >>
rect -25 24 -9 28
rect -25 -17 -21 24
rect -25 -21 -9 -17
<< ntransistor >>
rect -3 15 -1 21
<< ptransistor >>
rect -3 -13 -1 -7
<< polycontact >>
rect -5 8 -1 12
rect -5 -3 -1 1
<< ndcontact >>
rect -9 16 -5 20
rect 2 16 6 20
<< pdcontact >>
rect -9 -12 -5 -8
rect 2 -12 6 -8
<< m2contact >>
rect -9 24 -5 28
rect -9 -21 -5 -17
<< psubstratepcontact >>
rect -20 16 -16 20
<< nsubstratencontact >>
rect -18 -12 -14 -8
<< labels >>
rlabel metal1 -31 10 -31 10 3 A
rlabel metal1 -31 26 -31 26 4 in
rlabel metal1 12 6 12 6 7 out
rlabel metal1 -31 -10 -31 -10 3 vdd
rlabel metal1 -31 18 -31 18 3 gnd
rlabel metal1 -31 -1 -31 -1 3 Anot
<< end >>
