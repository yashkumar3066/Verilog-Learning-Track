magic
tech scmos
timestamp 1699384113
<< nwell >>
rect -7 16 58 37
<< polysilicon >>
rect 6 31 14 34
rect 36 31 44 34
rect 6 13 14 21
rect 6 8 7 13
rect 13 8 14 13
rect 6 -34 14 8
rect 36 -24 44 21
rect 36 -29 37 -24
rect 43 -29 44 -24
rect 36 -34 44 -29
rect 6 -46 14 -44
rect 36 -46 44 -44
<< ndiffusion >>
rect -4 -36 6 -34
rect -4 -42 -3 -36
rect 4 -42 6 -36
rect -4 -44 6 -42
rect 14 -36 36 -34
rect 14 -42 22 -36
rect 29 -42 36 -36
rect 14 -44 36 -42
rect 44 -36 55 -34
rect 44 -42 46 -36
rect 53 -42 55 -36
rect 44 -44 55 -42
<< pdiffusion >>
rect -4 29 6 31
rect -4 23 -3 29
rect 4 23 6 29
rect -4 21 6 23
rect 14 21 36 31
rect 44 29 55 31
rect 44 23 47 29
rect 54 23 55 29
rect 44 21 55 23
<< metal1 >>
rect -11 43 5 49
rect -4 29 5 43
rect -4 23 -3 29
rect 4 23 5 29
rect 46 29 55 30
rect 46 23 47 29
rect 54 23 55 29
rect -2 13 14 14
rect -2 8 7 13
rect 13 8 14 13
rect -2 7 14 8
rect 46 -1 55 23
rect 21 -10 60 -1
rect -3 -36 4 -35
rect -3 -52 4 -42
rect 21 -36 30 -10
rect 36 -24 53 -23
rect 36 -29 37 -24
rect 43 -29 53 -24
rect 36 -30 53 -29
rect 21 -42 22 -36
rect 29 -42 30 -36
rect 21 -43 30 -42
rect -9 -61 4 -52
<< ntransistor >>
rect 6 -44 14 -34
rect 36 -44 44 -34
<< ptransistor >>
rect 6 21 14 31
rect 36 21 44 31
<< polycontact >>
rect 7 8 13 13
rect 37 -29 43 -24
<< ndcontact >>
rect -3 -42 4 -36
rect 22 -42 29 -36
rect 46 -42 53 -36
<< pdcontact >>
rect -3 23 4 29
rect 47 23 54 29
<< labels >>
rlabel metal1 57 -6 57 -6 7 out
rlabel metal1 50 -27 50 -27 1 B
rlabel metal1 0 10 0 10 1 A
rlabel metal1 -6 -57 -6 -57 2 gnd
rlabel metal1 -4 45 -4 45 5 vdd
<< end >>
