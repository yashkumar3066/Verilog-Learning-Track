module \$_DLATCH_P_ (input E, input D, output Q);
  LATCH _TECHMAP_REPLACE_ (
  	.CLK(E),
  	.D(D),
  	.Q(Q)
  );
endmodule
